`timescale 1ns / 1ps

module rom (
    input  logic [31:0] addr,
    output logic [31:0] data
);
    logic [31:0] rom[0:15];

    initial begin
            rom[0] = 32'b00000000000000010100000010110111;
            rom[1] = 32'b00000000000000010100000010010111;
            rom[2] = 32'b00000001010000000000000011101111;
            rom[7] = 32'b00000000000000001000000011100111;
        // rom[0] = 32'b0000000_01000_00001_000_00100_0010011; //  r2 =8 + r1 
        // rom[1] = 32'b0000000_00100_11111_010_00100_0010011; //  r2 = 11 < r1 
        // rom[2] = 32'b0000000_01100_11111_011_00100_0010011; //  r2 =-signed < r1 
        // rom[3] = 32'b0000000_00100_00001_100_00100_0010011; //  r2 =8 ^ r1 
        // rom[4] = 32'b0000000_00111_00001_110_00100_0010011; //  r2 =8 | r1 
        // rom[5] = 32'b0000001_00000_00001_111_00100_0010011; //  r2 =8 & r1 
        // rom[6] = 32'b0000000_00001_00001_001_00100_0010011; //  r2 =r1 < 1
        // rom[7] = 32'b0000000_00001_00001_101_00100_0010011; //  r2 =r1 >> 1 
        // rom[8] = 32'b0100000_00011_00001_000_00100_0110011; //  r2 =r1 - r3 
        // rom[9] = 32'b0100000_00100_00010_101_00100_0010011; //  r2 =r1 >>> 4 

        // rom[0] = 32'b0000000_11111_00001_000_00001_0100011;
        // rom[1] = 32'b0000000_11111_00001_001_00001_0100011;
        // rom[2] = 32'b0000000_11111_00001_010_00001_0100011;
        // rom[3] = 32'b0000000_01100_00000_010_00100_0000011;
        // rom[4] = 32'b0000000_01100_00000_101_00100_0000011;
        //rtype
        // rom[1] = 32'b01000000001000001000001000110011;
        // rom[2] = 32'b00000000000111111010001000110011;
        // rom[3] = 32'b00000000000111111011001000110011;



        // rom[0] = 32'b00000000001000010000100001100011; // x6, x2, 8; x6 = 20
        // rom[4] = 32'b00000000001000010001100001100011;// x8 != x2, imm = 10 imode
        // rom[5] = 32'b00000000001111111100100001100011; // x8 != x2, imm = 10 imode
        // rom[9] = 32'b00000000001111111101100001100011; //bge x31, x3, 16
        // rom[10] = 32'b00000000001111111110100001100011; // x8 >= x2, imm = 10 imode
        // rom[11] = 32'b00000000001111111111100001100011; // x10 = x2-x8 
        // rom[15] = 32'b0000000_00010_01010_100_01000_1100011; // x10 < x2, imm = 10 imode
        // rom[17] = 32'b0000000_00010_01010_110_01000_1100011; // x10 < x2, imm = 10 imode unsinged

        
        // //rom[x]=32'b fucn7 _ rs2 _ rs1 _f3 _ rd  _opcode; // R-Type
        // rom[0] = 32'b0000000_00001_00010_000_00100_0110011; // add x4, x2, x1
        // rom[1] = 32'b0100000_00001_00010_000_00101_0110011; // sub x5, x2, x1
        // //rom[x]=32'b imm7  _ rs2 _ rs1 _f3 _ imm5_ opcode; // B-Type
        // rom[2] = 32'b0000000_00010_00010_000_01100_1100011; // beq x2, x2, 12 
        // //rom[x]=32'b imm7  _ rs2 _ rs1 _f3 _ imm5_ opcode; // S-Type
        // rom[3] = 32'b0000000_00010_00000_010_01000_0100011; // sw x2, 8(x0);
        // //rom[x]=32'b imm12      _ rs1 _f3 _ rd  _ opcode; // L-Type
        // rom[4] = 32'b000000001000_00000_010_00011_0000011; // lw x3, 8(x0);
        // //rom[x]=32'b imm12      _ rs1 _f3 _ rd  _ opcode; // I-Type
        // rom[5] = 32'b000000000001_00000_000_00001_0010011; // addi x1, x0, 1;
        // rom[6] = 32'b000000000010_00001_001_00110_0010011; // slli x6, x1, 2;
    end
    assign data = rom[addr[31:2]];
endmodule
